-- labmininios.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity labmininios is
	port (
		clk_clk         : in    std_logic                     := '0';             --       clk.clk
		h_bridge_export : out   std_logic_vector(2 downto 0);                     --  h_bridge.export
		lcd_export      : out   std_logic_vector(10 downto 0);                    --       lcd.export
		reset_reset     : in    std_logic                     := '0';             --     reset.reset
		sdram_addr      : out   std_logic_vector(12 downto 0);                    --     sdram.addr
		sdram_ba        : out   std_logic_vector(1 downto 0);                     --          .ba
		sdram_cas_n     : out   std_logic;                                        --          .cas_n
		sdram_cke       : out   std_logic;                                        --          .cke
		sdram_cs_n      : out   std_logic;                                        --          .cs_n
		sdram_dq        : inout std_logic_vector(15 downto 0) := (others => '0'); --          .dq
		sdram_dqm       : out   std_logic_vector(1 downto 0);                     --          .dqm
		sdram_ras_n     : out   std_logic;                                        --          .ras_n
		sdram_we_n      : out   std_logic;                                        --          .we_n
		sdram_clk_clk   : out   std_logic;                                        -- sdram_clk.clk
		switch_export   : in    std_logic_vector(9 downto 0)  := (others => '0')  --    switch.export
	);
end entity labmininios;

architecture rtl of labmininios is
	component labmininios_CPU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component labmininios_CPU;

	component labmininios_DMEM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component labmininios_DMEM;

	component labmininios_H_BRIDGE is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(2 downto 0)                      -- export
		);
	end component labmininios_H_BRIDGE;

	component labmininios_IMEM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component labmininios_IMEM;

	component labmininios_LCD is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(10 downto 0)                     -- export
		);
	end component labmininios_LCD;

	component labmininios_SWITCH is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component labmininios_SWITCH;

	component labmininios_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component labmininios_jtag_uart_0;

	component labmininios_sys_sdram_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component labmininios_sys_sdram_pll_0;

	component labmininios_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component labmininios_sysid_qsys_0;

	component labmininios_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component labmininios_timer_0;

	component labmininios_mm_interconnect_0 is
		port (
			sys_sdram_pll_0_sys_clk_clk               : in  std_logic                     := 'X';             -- clk
			CPU_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			CPU_data_master_address                   : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			CPU_data_master_waitrequest               : out std_logic;                                        -- waitrequest
			CPU_data_master_byteenable                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_master_read                      : in  std_logic                     := 'X';             -- read
			CPU_data_master_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_master_write                     : in  std_logic                     := 'X';             -- write
			CPU_data_master_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_master_debugaccess               : in  std_logic                     := 'X';             -- debugaccess
			CPU_instruction_master_address            : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			CPU_instruction_master_waitrequest        : out std_logic;                                        -- waitrequest
			CPU_instruction_master_read               : in  std_logic                     := 'X';             -- read
			CPU_instruction_master_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_debug_mem_slave_address               : out std_logic_vector(8 downto 0);                     -- address
			CPU_debug_mem_slave_write                 : out std_logic;                                        -- write
			CPU_debug_mem_slave_read                  : out std_logic;                                        -- read
			CPU_debug_mem_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_debug_mem_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_debug_mem_slave_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_debug_mem_slave_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			CPU_debug_mem_slave_debugaccess           : out std_logic;                                        -- debugaccess
			DMEM_s1_address                           : out std_logic_vector(24 downto 0);                    -- address
			DMEM_s1_write                             : out std_logic;                                        -- write
			DMEM_s1_read                              : out std_logic;                                        -- read
			DMEM_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			DMEM_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			DMEM_s1_byteenable                        : out std_logic_vector(1 downto 0);                     -- byteenable
			DMEM_s1_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			DMEM_s1_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			DMEM_s1_chipselect                        : out std_logic;                                        -- chipselect
			H_BRIDGE_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			H_BRIDGE_s1_write                         : out std_logic;                                        -- write
			H_BRIDGE_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			H_BRIDGE_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			H_BRIDGE_s1_chipselect                    : out std_logic;                                        -- chipselect
			IMEM_s1_address                           : out std_logic_vector(15 downto 0);                    -- address
			IMEM_s1_write                             : out std_logic;                                        -- write
			IMEM_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			IMEM_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			IMEM_s1_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			IMEM_s1_chipselect                        : out std_logic;                                        -- chipselect
			IMEM_s1_clken                             : out std_logic;                                        -- clken
			jtag_uart_0_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			LCD_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			LCD_s1_write                              : out std_logic;                                        -- write
			LCD_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LCD_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			LCD_s1_chipselect                         : out std_logic;                                        -- chipselect
			SWITCH_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			SWITCH_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_qsys_0_control_slave_address        : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                        : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                          : out std_logic;                                        -- write
			timer_0_s1_readdata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                      : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                     : out std_logic                                         -- chipselect
		);
	end component labmininios_mm_interconnect_0;

	component labmininios_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component labmininios_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal sys_sdram_pll_0_sys_clk_clk                                     : std_logic;                     -- sys_sdram_pll_0:sys_clk_clk -> [CPU:clk, DMEM:clk, H_BRIDGE:clk, IMEM:clk, LCD:clk, SWITCH:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, rst_controller:clk, sysid_qsys_0:clock, timer_0:clk]
	signal cpu_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	signal cpu_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_debugaccess                                     : std_logic;                     -- CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	signal cpu_data_master_address                                         : std_logic_vector(26 downto 0); -- CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	signal cpu_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	signal cpu_data_master_read                                            : std_logic;                     -- CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	signal cpu_data_master_write                                           : std_logic;                     -- CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	signal cpu_data_master_writedata                                       : std_logic_vector(31 downto 0); -- CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	signal cpu_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	signal cpu_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                  : std_logic_vector(26 downto 0); -- CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	signal cpu_instruction_master_read                                     : std_logic;                     -- CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest               : std_logic;                     -- CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	signal mm_interconnect_0_imem_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:IMEM_s1_chipselect -> IMEM:chipselect
	signal mm_interconnect_0_imem_s1_readdata                              : std_logic_vector(31 downto 0); -- IMEM:readdata -> mm_interconnect_0:IMEM_s1_readdata
	signal mm_interconnect_0_imem_s1_address                               : std_logic_vector(15 downto 0); -- mm_interconnect_0:IMEM_s1_address -> IMEM:address
	signal mm_interconnect_0_imem_s1_byteenable                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:IMEM_s1_byteenable -> IMEM:byteenable
	signal mm_interconnect_0_imem_s1_write                                 : std_logic;                     -- mm_interconnect_0:IMEM_s1_write -> IMEM:write
	signal mm_interconnect_0_imem_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:IMEM_s1_writedata -> IMEM:writedata
	signal mm_interconnect_0_imem_s1_clken                                 : std_logic;                     -- mm_interconnect_0:IMEM_s1_clken -> IMEM:clken
	signal mm_interconnect_0_dmem_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:DMEM_s1_chipselect -> DMEM:az_cs
	signal mm_interconnect_0_dmem_s1_readdata                              : std_logic_vector(15 downto 0); -- DMEM:za_data -> mm_interconnect_0:DMEM_s1_readdata
	signal mm_interconnect_0_dmem_s1_waitrequest                           : std_logic;                     -- DMEM:za_waitrequest -> mm_interconnect_0:DMEM_s1_waitrequest
	signal mm_interconnect_0_dmem_s1_address                               : std_logic_vector(24 downto 0); -- mm_interconnect_0:DMEM_s1_address -> DMEM:az_addr
	signal mm_interconnect_0_dmem_s1_read                                  : std_logic;                     -- mm_interconnect_0:DMEM_s1_read -> mm_interconnect_0_dmem_s1_read:in
	signal mm_interconnect_0_dmem_s1_byteenable                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:DMEM_s1_byteenable -> mm_interconnect_0_dmem_s1_byteenable:in
	signal mm_interconnect_0_dmem_s1_readdatavalid                         : std_logic;                     -- DMEM:za_valid -> mm_interconnect_0:DMEM_s1_readdatavalid
	signal mm_interconnect_0_dmem_s1_write                                 : std_logic;                     -- mm_interconnect_0:DMEM_s1_write -> mm_interconnect_0_dmem_s1_write:in
	signal mm_interconnect_0_dmem_s1_writedata                             : std_logic_vector(15 downto 0); -- mm_interconnect_0:DMEM_s1_writedata -> DMEM:az_data
	signal mm_interconnect_0_timer_0_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                           : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                              : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_h_bridge_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:H_BRIDGE_s1_chipselect -> H_BRIDGE:chipselect
	signal mm_interconnect_0_h_bridge_s1_readdata                          : std_logic_vector(31 downto 0); -- H_BRIDGE:readdata -> mm_interconnect_0:H_BRIDGE_s1_readdata
	signal mm_interconnect_0_h_bridge_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:H_BRIDGE_s1_address -> H_BRIDGE:address
	signal mm_interconnect_0_h_bridge_s1_write                             : std_logic;                     -- mm_interconnect_0:H_BRIDGE_s1_write -> mm_interconnect_0_h_bridge_s1_write:in
	signal mm_interconnect_0_h_bridge_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:H_BRIDGE_s1_writedata -> H_BRIDGE:writedata
	signal mm_interconnect_0_lcd_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:LCD_s1_chipselect -> LCD:chipselect
	signal mm_interconnect_0_lcd_s1_readdata                               : std_logic_vector(31 downto 0); -- LCD:readdata -> mm_interconnect_0:LCD_s1_readdata
	signal mm_interconnect_0_lcd_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LCD_s1_address -> LCD:address
	signal mm_interconnect_0_lcd_s1_write                                  : std_logic;                     -- mm_interconnect_0:LCD_s1_write -> mm_interconnect_0_lcd_s1_write:in
	signal mm_interconnect_0_lcd_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:LCD_s1_writedata -> LCD:writedata
	signal mm_interconnect_0_switch_s1_readdata                            : std_logic_vector(31 downto 0); -- SWITCH:readdata -> mm_interconnect_0:SWITCH_s1_readdata
	signal mm_interconnect_0_switch_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SWITCH_s1_address -> SWITCH:address
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- timer_0:irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [IMEM:reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [CPU:reset_req, IMEM:reset_req, rst_translator:reset_req_in]
	signal sys_sdram_pll_0_reset_source_reset                              : std_logic;                     -- sys_sdram_pll_0:reset_source_reset -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_dmem_s1_read_ports_inv                        : std_logic;                     -- mm_interconnect_0_dmem_s1_read:inv -> DMEM:az_rd_n
	signal mm_interconnect_0_dmem_s1_byteenable_ports_inv                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0_dmem_s1_byteenable:inv -> DMEM:az_be_n
	signal mm_interconnect_0_dmem_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_dmem_s1_write:inv -> DMEM:az_wr_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_h_bridge_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_h_bridge_s1_write:inv -> H_BRIDGE:write_n
	signal mm_interconnect_0_lcd_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_lcd_s1_write:inv -> LCD:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [CPU:reset_n, DMEM:reset_n, H_BRIDGE:reset_n, LCD:reset_n, SWITCH:reset_n, jtag_uart_0:rst_n, sysid_qsys_0:reset_n, timer_0:reset_n]

begin

	cpu : component labmininios_CPU
		port map (
			clk                                 => sys_sdram_pll_0_sys_clk_clk,                       --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                              --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	dmem : component labmininios_DMEM
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                    --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,       -- reset.reset_n
			az_addr        => mm_interconnect_0_dmem_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_dmem_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_dmem_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_dmem_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_dmem_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_dmem_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_dmem_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_dmem_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_dmem_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                     --  wire.export
			zs_ba          => sdram_ba,                                       --      .export
			zs_cas_n       => sdram_cas_n,                                    --      .export
			zs_cke         => sdram_cke,                                      --      .export
			zs_cs_n        => sdram_cs_n,                                     --      .export
			zs_dq          => sdram_dq,                                       --      .export
			zs_dqm         => sdram_dqm,                                      --      .export
			zs_ras_n       => sdram_ras_n,                                    --      .export
			zs_we_n        => sdram_we_n                                      --      .export
		);

	h_bridge : component labmininios_H_BRIDGE
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_h_bridge_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_h_bridge_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_h_bridge_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_h_bridge_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_h_bridge_s1_readdata,        --                    .readdata
			out_port   => h_bridge_export                                -- external_connection.export
		);

	imem : component labmininios_IMEM
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,          --   clk1.clk
			address    => mm_interconnect_0_imem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_imem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_imem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_imem_s1_write,      --       .write
			readdata   => mm_interconnect_0_imem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_imem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_imem_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,       -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,   --       .reset_req
			freeze     => '0'                                   -- (terminated)
		);

	lcd : component labmininios_LCD
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_lcd_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_lcd_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_lcd_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_lcd_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_lcd_s1_readdata,        --                    .readdata
			out_port   => lcd_export                                -- external_connection.export
		);

	switch : component labmininios_SWITCH
		port map (
			clk      => sys_sdram_pll_0_sys_clk_clk,              --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switch_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_switch_s1_readdata,     --                    .readdata
			in_port  => switch_export                             -- external_connection.export
		);

	jtag_uart_0 : component labmininios_jtag_uart_0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                     --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	sys_sdram_pll_0 : component labmininios_sys_sdram_pll_0
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => reset_reset,                        --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                      --    sdram_clk.clk
			reset_source_reset => sys_sdram_pll_0_reset_source_reset  -- reset_source.reset
		);

	sysid_qsys_0 : component labmininios_sysid_qsys_0
		port map (
			clock    => sys_sdram_pll_0_sys_clk_clk,                             --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	timer_0 : component labmininios_timer_0
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                  --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	mm_interconnect_0 : component labmininios_mm_interconnect_0
		port map (
			sys_sdram_pll_0_sys_clk_clk               => sys_sdram_pll_0_sys_clk_clk,                                 --         sys_sdram_pll_0_sys_clk.clk
			CPU_reset_reset_bridge_in_reset_reset     => rst_controller_reset_out_reset,                              -- CPU_reset_reset_bridge_in_reset.reset
			CPU_data_master_address                   => cpu_data_master_address,                                     --                 CPU_data_master.address
			CPU_data_master_waitrequest               => cpu_data_master_waitrequest,                                 --                                .waitrequest
			CPU_data_master_byteenable                => cpu_data_master_byteenable,                                  --                                .byteenable
			CPU_data_master_read                      => cpu_data_master_read,                                        --                                .read
			CPU_data_master_readdata                  => cpu_data_master_readdata,                                    --                                .readdata
			CPU_data_master_write                     => cpu_data_master_write,                                       --                                .write
			CPU_data_master_writedata                 => cpu_data_master_writedata,                                   --                                .writedata
			CPU_data_master_debugaccess               => cpu_data_master_debugaccess,                                 --                                .debugaccess
			CPU_instruction_master_address            => cpu_instruction_master_address,                              --          CPU_instruction_master.address
			CPU_instruction_master_waitrequest        => cpu_instruction_master_waitrequest,                          --                                .waitrequest
			CPU_instruction_master_read               => cpu_instruction_master_read,                                 --                                .read
			CPU_instruction_master_readdata           => cpu_instruction_master_readdata,                             --                                .readdata
			CPU_debug_mem_slave_address               => mm_interconnect_0_cpu_debug_mem_slave_address,               --             CPU_debug_mem_slave.address
			CPU_debug_mem_slave_write                 => mm_interconnect_0_cpu_debug_mem_slave_write,                 --                                .write
			CPU_debug_mem_slave_read                  => mm_interconnect_0_cpu_debug_mem_slave_read,                  --                                .read
			CPU_debug_mem_slave_readdata              => mm_interconnect_0_cpu_debug_mem_slave_readdata,              --                                .readdata
			CPU_debug_mem_slave_writedata             => mm_interconnect_0_cpu_debug_mem_slave_writedata,             --                                .writedata
			CPU_debug_mem_slave_byteenable            => mm_interconnect_0_cpu_debug_mem_slave_byteenable,            --                                .byteenable
			CPU_debug_mem_slave_waitrequest           => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,           --                                .waitrequest
			CPU_debug_mem_slave_debugaccess           => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,           --                                .debugaccess
			DMEM_s1_address                           => mm_interconnect_0_dmem_s1_address,                           --                         DMEM_s1.address
			DMEM_s1_write                             => mm_interconnect_0_dmem_s1_write,                             --                                .write
			DMEM_s1_read                              => mm_interconnect_0_dmem_s1_read,                              --                                .read
			DMEM_s1_readdata                          => mm_interconnect_0_dmem_s1_readdata,                          --                                .readdata
			DMEM_s1_writedata                         => mm_interconnect_0_dmem_s1_writedata,                         --                                .writedata
			DMEM_s1_byteenable                        => mm_interconnect_0_dmem_s1_byteenable,                        --                                .byteenable
			DMEM_s1_readdatavalid                     => mm_interconnect_0_dmem_s1_readdatavalid,                     --                                .readdatavalid
			DMEM_s1_waitrequest                       => mm_interconnect_0_dmem_s1_waitrequest,                       --                                .waitrequest
			DMEM_s1_chipselect                        => mm_interconnect_0_dmem_s1_chipselect,                        --                                .chipselect
			H_BRIDGE_s1_address                       => mm_interconnect_0_h_bridge_s1_address,                       --                     H_BRIDGE_s1.address
			H_BRIDGE_s1_write                         => mm_interconnect_0_h_bridge_s1_write,                         --                                .write
			H_BRIDGE_s1_readdata                      => mm_interconnect_0_h_bridge_s1_readdata,                      --                                .readdata
			H_BRIDGE_s1_writedata                     => mm_interconnect_0_h_bridge_s1_writedata,                     --                                .writedata
			H_BRIDGE_s1_chipselect                    => mm_interconnect_0_h_bridge_s1_chipselect,                    --                                .chipselect
			IMEM_s1_address                           => mm_interconnect_0_imem_s1_address,                           --                         IMEM_s1.address
			IMEM_s1_write                             => mm_interconnect_0_imem_s1_write,                             --                                .write
			IMEM_s1_readdata                          => mm_interconnect_0_imem_s1_readdata,                          --                                .readdata
			IMEM_s1_writedata                         => mm_interconnect_0_imem_s1_writedata,                         --                                .writedata
			IMEM_s1_byteenable                        => mm_interconnect_0_imem_s1_byteenable,                        --                                .byteenable
			IMEM_s1_chipselect                        => mm_interconnect_0_imem_s1_chipselect,                        --                                .chipselect
			IMEM_s1_clken                             => mm_interconnect_0_imem_s1_clken,                             --                                .clken
			jtag_uart_0_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --   jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                .write
			jtag_uart_0_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                .read
			jtag_uart_0_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                .readdata
			jtag_uart_0_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                .chipselect
			LCD_s1_address                            => mm_interconnect_0_lcd_s1_address,                            --                          LCD_s1.address
			LCD_s1_write                              => mm_interconnect_0_lcd_s1_write,                              --                                .write
			LCD_s1_readdata                           => mm_interconnect_0_lcd_s1_readdata,                           --                                .readdata
			LCD_s1_writedata                          => mm_interconnect_0_lcd_s1_writedata,                          --                                .writedata
			LCD_s1_chipselect                         => mm_interconnect_0_lcd_s1_chipselect,                         --                                .chipselect
			SWITCH_s1_address                         => mm_interconnect_0_switch_s1_address,                         --                       SWITCH_s1.address
			SWITCH_s1_readdata                        => mm_interconnect_0_switch_s1_readdata,                        --                                .readdata
			sysid_qsys_0_control_slave_address        => mm_interconnect_0_sysid_qsys_0_control_slave_address,        --      sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata       => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,       --                                .readdata
			timer_0_s1_address                        => mm_interconnect_0_timer_0_s1_address,                        --                      timer_0_s1.address
			timer_0_s1_write                          => mm_interconnect_0_timer_0_s1_write,                          --                                .write
			timer_0_s1_readdata                       => mm_interconnect_0_timer_0_s1_readdata,                       --                                .readdata
			timer_0_s1_writedata                      => mm_interconnect_0_timer_0_s1_writedata,                      --                                .writedata
			timer_0_s1_chipselect                     => mm_interconnect_0_timer_0_s1_chipselect                      --                                .chipselect
		);

	irq_mapper : component labmininios_irq_mapper
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,    --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_sdram_pll_0_reset_source_reset, -- reset_in0.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_dmem_s1_read_ports_inv <= not mm_interconnect_0_dmem_s1_read;

	mm_interconnect_0_dmem_s1_byteenable_ports_inv <= not mm_interconnect_0_dmem_s1_byteenable;

	mm_interconnect_0_dmem_s1_write_ports_inv <= not mm_interconnect_0_dmem_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_h_bridge_s1_write_ports_inv <= not mm_interconnect_0_h_bridge_s1_write;

	mm_interconnect_0_lcd_s1_write_ports_inv <= not mm_interconnect_0_lcd_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of labmininios
